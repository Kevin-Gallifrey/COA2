`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/04/23 15:09:16
// Design Name: 
// Module Name: CU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module CU(
    input clk,
    input rst,
    input [7:0] IR,
    output  [16:0] C,
    output  [3:0] OP
    );
    
    //  control memory
    reg [20:0] CM [0:92];
    //CM[][20:17]=Op[3:0] CM[][16:0]=C16~C0
    
	parameter idle=0, decode=1, fetch=2, run=3;
	reg [1:0] step=0;
	reg [7:0] CAR=0;
	reg [20:0] CBR=0;
    
    parameter STORE_X=1, LOAD_X=2;
    
      assign OP = CBR[20:17];
     assign C = CBR[16:0];
     
    always@(posedge clk or negedge rst)
	begin
        if(~rst)
            begin
                step <= idle;
                //��ʼ��CM
                //Fetch Instruction
                CM[0]=21'b000000000010000000001;
                CM[1]=21'b000000000000000001001;
                CM[2]=21'b000000000000000010001;
                CM[3]=21'b000000000000001000010;
                //STORE X
                CM[4]=21'b000000000000000100001;
                CM[5]=21'b000000000100000000001;
                CM[6]=21'b000000001000000000100;
                //LOAD [X]
                CM[7]=21'b000000000000000100001;
                CM[8]=21'b000000000000000001001;
                CM[9]=21'b000000000000110000001;
                CM[10]=21'b011001100000000000001;
                CM[11]=21'b000010000000000000100;
                //ADD [X]
                CM[12]=21'b000000000000000100001;
                CM[13]=21'b000000000000000001001;
                CM[14]=21'b000000000000010000001;
                CM[15]=21'b000101100000000000001;
                CM[16]=21'b000010000000000000100;
                //SUB [X]
                CM[17]=21'b000000000000000100001;
                CM[18]=21'b000000000000000001001;
                CM[19]=21'b000000000000010000001;
                CM[20]=21'b001001100000000000001;
                CM[21]=21'b000010000000000000100;
                //JMPGEZ X(ACC<0)
                CM[22]=21'b000000000000000000100;
                //JMP X & JMPGEZ X(ACC��0)
                CM[23]=21'b000000010000000000100;
                //HALT
                CM[24]=21'b000000000000000000000;
                //MPY [X]
                CM[25]=21'b000000000000000100001;
                CM[26]=21'b000000000000000001001;
                CM[27]=21'b000000000000010000001;
                CM[28]=21'b001101100000000000001;
                CM[29]=21'b000010000000000000100;
                //DIV [X]
                CM[30]=21'b000000000000000100001;
                CM[31]=21'b000000000000000001001;
                CM[32]=21'b000000000000010000001;
                CM[33]=21'b010001100000000000001;
                CM[34]=21'b000010000000000000100;
                //AND [X]
                CM[35]=21'b000000000000000100001;
                CM[36]=21'b000000000000000001001;
                CM[37]=21'b000000000000010000001;
                CM[38]=21'b010101100000000000001;
                CM[39]=21'b000010000000000000100;
                //OR [X]
                CM[40]=21'b000000000000000100001;
                CM[41]=21'b000000000000000001001;
                CM[42]=21'b000000000000010000001;
                CM[43]=21'b011001100000000000001;
                CM[44]=21'b000010000000000000100;
                //XOR [X]
                CM[45]=21'b000000000000000100001;
                CM[46]=21'b000000000000000001001;
                CM[47]=21'b000000000000010000001;
                CM[48]=21'b011101100000000000001;
                CM[49]=21'b000010000000000000100;
                //NOT [X]
                CM[50]=21'b000000000000000100001;
                CM[51]=21'b000000000000000001001;
                CM[52]=21'b000000000000010000001;
                CM[53]=21'b100000100000000000001;
                CM[54]=21'b000010000000000000100;
                //SHIFTR
                CM[55]=21'b100101000000000000100;
                //SHIFTL
                CM[56]=21'b101001000000000000100;
                //LOAD X
                CM[57]=21'b000000000000110000001;
                CM[58]=21'b000000000001000000001;
                CM[59]=21'b011001100000000000001;
                CM[60]=21'b000010000000000000100;
                //ADD X
                CM[61]=21'b000000000000010000001;
                CM[62]=21'b000000000001000000001;
                CM[63]=21'b000101100000000000001;
                CM[64]=21'b000010000000000000100;
                //SUB X
                CM[65]=21'b000000000000010000001;
                CM[66]=21'b000000000001000000001;
                CM[67]=21'b001001100000000000001;
                CM[68]=21'b000010000000000000100;
                //MPY X
                CM[69]=21'b000000000000010000001;
                CM[70]=21'b000000000001000000001;
                CM[71]=21'b001101100000000000001;
                CM[72]=21'b000010000000000000100;
                //DIV X
                CM[73]=21'b000000000000010000001;
                CM[74]=21'b000000000001000000001;
                CM[75]=21'b010001100000000000001;
                CM[76]=21'b000010000000000000100;
                //AND X
                CM[77]=21'b000000000000010000001;
                CM[78]=21'b000000000001000000001;
                CM[79]=21'b010101100000000000001;
                CM[80]=21'b000010000000000000100;
                //OR X
                CM[81]=21'b000000000000010000001;
                CM[82]=21'b000000000001000000001;
                CM[83]=21'b011001100000000000001;
                CM[84]=21'b000010000000000000100;
                //XOR X
                CM[85]=21'b000000000000010000001;
                CM[86]=21'b000000000001000000001;
                CM[87]=21'b011101100000000000001;
                CM[88]=21'b000010000000000000100;
                //NOT X
                CM[89]=21'b000000000000010000001;
                CM[90]=21'b000000000001000000001;
                CM[91]=21'b100001100000000000001;
                CM[92]=21'b000010000000000000100;
            end
        else
        begin
            case(step)
                idle:begin
                    CAR <= 0;
                    CBR <= 0;
                    step <= fetch;
                end
                //���룬��IR�õ�CM��΢ָ��ĵ�ַ?
                decode:begin
                    case(IR)
                        STORE_X:begin
                        $display("STORE X");
                            CAR <= 4;
                            step <= fetch;
                        end
                        LOAD_X:begin
                         $display("LOAD X");
                            CAR <= 7;
                            step <= fetch;
                        end                        
                        default: step <= idle;	//û����Чָ�����idle
                    endcase
                end
                //ȡָ�����CARȡ��΢ָ�CBR
                fetch:begin
                    CBR <= CM[CAR];
                    step <= run;
                end
                //����΢ָ���������źŲ��õ���һ��΢ָ��ĵ�ַ?
                run:begin
                    CBR <= 0;
                    case(CBR[2:0])
                        3'b001:begin
                            CAR <= CAR + 1;
                            step <= fetch;
                        end
                        3'b010:begin
                            step <= decode;
                        end
                        3'b100:begin
                            CAR <= 0;
                            step <= fetch;
                        end
                        default:begin
                            step <= idle;
                        end
                    endcase
                end
                
            endcase
        end
    end
	
endmodule